`ifndef IMPORTED_CLN_TXC_STRUCTS
`define IMPORTED_CLN_TXC_STRUCTS
import CLN_TXC_structs::*;
`endif
