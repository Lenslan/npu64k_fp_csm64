
module npu_tb_top();
    core_chip_tb u_core_chip_tb();

endmodule: npu_tb_top
