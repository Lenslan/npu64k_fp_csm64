`ifndef IMPORTED_CLN_STRUCTS
`define IMPORTED_CLN_STRUCTS
import CLN_structs::*;
`endif
